// A simple ALU

module day4 (
	input     logic [7:0]   a_i,
	input     logic [7:0]   b_i,
	input     logic [2:0]   op_i,

	output    logic [7:0]   alu_o
);

	// Write your logic here...

endmodule
