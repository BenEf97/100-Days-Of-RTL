// Simple ALU TB

module day4_tb ();

  // Write your Testbench here...

endmodule
